module mnist_classifier (
    input wire clk,
    input wire rst_n,
    input wire start,              
    output reg [9:0] ram_addr,     
    input wire       ram_data,     
    output reg [3:0] prediction,   
    output reg       done          
);

    localparam IDLE = 0, WAIT_RAM = 1, CALC = 2, RESULT = 3;
    reg [1:0] state;
    
    reg signed [15:0] score [0:9];
    reg [9:0] total_ink;

    reg [9:0] rom_data;         
    reg [9:0] rom_data_left;    
    reg [9:0] rom_data_right;   
    
    // --- FUNÇÃO CORRIGIDA (SINTAXE ROBUSTA) ---
    function [9:0] get_rom_data;
        input [9:0] addr;
        begin
        case (addr)
            10'd0   : rom_data = 10'b0000000000;
            10'd1   : rom_data = 10'b0000000000;
            10'd2   : rom_data = 10'b0000000000;
            10'd3   : rom_data = 10'b0000000000;
            10'd4   : rom_data = 10'b0000000000;
            10'd5   : rom_data = 10'b0000000000;
            10'd6   : rom_data = 10'b0000000000;
            10'd7   : rom_data = 10'b0000000000;
            10'd8   : rom_data = 10'b0000000000;
            10'd9   : rom_data = 10'b0000000000;
            10'd10  : rom_data = 10'b0000000000;
            10'd11  : rom_data = 10'b0000000000;
            10'd12  : rom_data = 10'b0000000000;
            10'd13  : rom_data = 10'b0000000000;
            10'd14  : rom_data = 10'b0000000000;
            10'd15  : rom_data = 10'b0000000000;
            10'd16  : rom_data = 10'b0000000000;
            10'd17  : rom_data = 10'b0000000000;
            10'd18  : rom_data = 10'b0000000000;
            10'd19  : rom_data = 10'b0000000000;
            10'd20  : rom_data = 10'b0000000000;
            10'd21  : rom_data = 10'b0000000000;
            10'd22  : rom_data = 10'b0000000000;
            10'd23  : rom_data = 10'b0000000000;
            10'd24  : rom_data = 10'b0000000000;
            10'd25  : rom_data = 10'b0000000000;
            10'd26  : rom_data = 10'b0000000000;
            10'd27  : rom_data = 10'b0000000000;
            10'd28  : rom_data = 10'b0000000000;
            10'd29  : rom_data = 10'b0000000000;
            10'd30  : rom_data = 10'b0000000000;
            10'd31  : rom_data = 10'b0000000000;
            10'd32  : rom_data = 10'b0000000000;
            10'd33  : rom_data = 10'b0000000000;
            10'd34  : rom_data = 10'b0000000000;
            10'd35  : rom_data = 10'b0000000000;
            10'd36  : rom_data = 10'b0000000000;
            10'd37  : rom_data = 10'b0000000000;
            10'd38  : rom_data = 10'b0000000000;
            10'd39  : rom_data = 10'b0000000000;
            10'd40  : rom_data = 10'b0000000000;
            10'd41  : rom_data = 10'b0000000000;
            10'd42  : rom_data = 10'b0000000000;
            10'd43  : rom_data = 10'b0000000000;
            10'd44  : rom_data = 10'b0000000000;
            10'd45  : rom_data = 10'b0000000000;
            10'd46  : rom_data = 10'b0000000000;
            10'd47  : rom_data = 10'b0000000000;
            10'd48  : rom_data = 10'b0000000000;
            10'd49  : rom_data = 10'b0000000000;
            10'd50  : rom_data = 10'b0000000000;
            10'd51  : rom_data = 10'b0000000000;
            10'd52  : rom_data = 10'b0000000000;
            10'd53  : rom_data = 10'b0000000000;
            10'd54  : rom_data = 10'b0000000000;
            10'd55  : rom_data = 10'b0000000000;
            10'd56  : rom_data = 10'b0000000000;
            10'd57  : rom_data = 10'b0000000000;
            10'd58  : rom_data = 10'b0000000000;
            10'd59  : rom_data = 10'b0000000000;
            10'd60  : rom_data = 10'b0000000000;
            10'd61  : rom_data = 10'b0000000000;
            10'd62  : rom_data = 10'b0000000000;
            10'd63  : rom_data = 10'b0000000000;
            10'd64  : rom_data = 10'b0000000000;
            10'd65  : rom_data = 10'b0000000000;
            10'd66  : rom_data = 10'b0000000000;
            10'd67  : rom_data = 10'b0000000000;
            10'd68  : rom_data = 10'b0000000000;
            10'd69  : rom_data = 10'b0000000000;
            10'd70  : rom_data = 10'b0000000000;
            10'd71  : rom_data = 10'b0000000000;
            10'd72  : rom_data = 10'b0000000000;
            10'd73  : rom_data = 10'b0000000000;
            10'd74  : rom_data = 10'b0000000000;
            10'd75  : rom_data = 10'b0000000000;
            10'd76  : rom_data = 10'b0000000000;
            10'd77  : rom_data = 10'b0000000000;
            10'd78  : rom_data = 10'b0000000000;
            10'd79  : rom_data = 10'b0000000000;
            10'd80  : rom_data = 10'b0000000000;
            10'd81  : rom_data = 10'b0000000000;
            10'd82  : rom_data = 10'b0000000000;
            10'd83  : rom_data = 10'b0000000000;
            10'd84  : rom_data = 10'b0000000000;
            10'd85  : rom_data = 10'b0000000000;
            10'd86  : rom_data = 10'b0000000000;
            10'd87  : rom_data = 10'b0000000000;
            10'd88  : rom_data = 10'b0000000000;
            10'd89  : rom_data = 10'b0000000000;
            10'd90  : rom_data = 10'b0000000000;
            10'd91  : rom_data = 10'b0000000000;
            10'd92  : rom_data = 10'b0000000000;
            10'd93  : rom_data = 10'b0000000000;
            10'd94  : rom_data = 10'b0000000000;
            10'd95  : rom_data = 10'b0000000000;
            10'd96  : rom_data = 10'b0000000000;
            10'd97  : rom_data = 10'b0000000000;
            10'd98  : rom_data = 10'b0000000000;
            10'd99  : rom_data = 10'b0000000000;
            10'd100 : rom_data = 10'b0000000000;
            10'd101 : rom_data = 10'b0000000000;
            10'd102 : rom_data = 10'b0000000000;
            10'd103 : rom_data = 10'b0000000000;
            10'd104 : rom_data = 10'b0000000000;
            10'd105 : rom_data = 10'b0000000000;
            10'd106 : rom_data = 10'b0000000000;
            10'd107 : rom_data = 10'b0000000000;
            10'd108 : rom_data = 10'b0000000000;
            10'd109 : rom_data = 10'b0000000000;
            10'd110 : rom_data = 10'b0000000000;
            10'd111 : rom_data = 10'b0000000000;
            10'd112 : rom_data = 10'b0000000000;
            10'd113 : rom_data = 10'b0000000000;
            10'd114 : rom_data = 10'b0000000000;
            10'd115 : rom_data = 10'b0000000000;
            10'd116 : rom_data = 10'b0000000000;
            10'd117 : rom_data = 10'b0000000000;
            10'd118 : rom_data = 10'b0000000000;
            10'd119 : rom_data = 10'b0000000000;
            10'd120 : rom_data = 10'b0000000000;
            10'd121 : rom_data = 10'b0000000000;
            10'd122 : rom_data = 10'b0000000000;
            10'd123 : rom_data = 10'b0000000000;
            10'd124 : rom_data = 10'b0000000100;
            10'd125 : rom_data = 10'b0000000100;
            10'd126 : rom_data = 10'b0001000100;
            10'd127 : rom_data = 10'b0001000100;
            10'd128 : rom_data = 10'b0001000100;
            10'd129 : rom_data = 10'b0001000100;
            10'd130 : rom_data = 10'b0000000000;
            10'd131 : rom_data = 10'b0000000000;
            10'd132 : rom_data = 10'b0000000000;
            10'd133 : rom_data = 10'b0000000000;
            10'd134 : rom_data = 10'b0000000000;
            10'd135 : rom_data = 10'b0000000000;
            10'd136 : rom_data = 10'b0000000000;
            10'd137 : rom_data = 10'b0000000000;
            10'd138 : rom_data = 10'b0000000000;
            10'd139 : rom_data = 10'b0000000000;
            10'd140 : rom_data = 10'b0000000000;
            10'd141 : rom_data = 10'b0000000000;
            10'd142 : rom_data = 10'b0000000000;
            10'd143 : rom_data = 10'b0000000000;
            10'd144 : rom_data = 10'b0000000000;
            10'd145 : rom_data = 10'b0000000000;
            10'd146 : rom_data = 10'b0000000000;
            10'd147 : rom_data = 10'b0000000000;
            10'd148 : rom_data = 10'b0000000000;
            10'd149 : rom_data = 10'b0000000000;
            10'd150 : rom_data = 10'b0000001100;
            10'd151 : rom_data = 10'b0000001100;
            10'd152 : rom_data = 10'b0000001100;
            10'd153 : rom_data = 10'b0101001101;
            10'd154 : rom_data = 10'b0101001101;
            10'd155 : rom_data = 10'b0101001111;
            10'd156 : rom_data = 10'b0101001111;
            10'd157 : rom_data = 10'b0101001101;
            10'd158 : rom_data = 10'b0100000101;
            10'd159 : rom_data = 10'b0000000001;
            10'd160 : rom_data = 10'b0000000000;
            10'd161 : rom_data = 10'b0000000000;
            10'd162 : rom_data = 10'b0000000000;
            10'd163 : rom_data = 10'b0000000000;
            10'd164 : rom_data = 10'b0000000000;
            10'd165 : rom_data = 10'b0000000000;
            10'd166 : rom_data = 10'b0000000000;
            10'd167 : rom_data = 10'b0000000000;
            10'd168 : rom_data = 10'b0000000000;
            10'd169 : rom_data = 10'b0000000000;
            10'd170 : rom_data = 10'b0000000000;
            10'd171 : rom_data = 10'b0000000000;
            10'd172 : rom_data = 10'b0000000000;
            10'd173 : rom_data = 10'b0000000000;
            10'd174 : rom_data = 10'b0000000000;
            10'd175 : rom_data = 10'b0000000000;
            10'd176 : rom_data = 10'b0000000000;
            10'd177 : rom_data = 10'b0000001100;
            10'd178 : rom_data = 10'b0000001100;
            10'd179 : rom_data = 10'b0100001100;
            10'd180 : rom_data = 10'b0101101101;
            10'd181 : rom_data = 10'b0101101101;
            10'd182 : rom_data = 10'b1101101111;
            10'd183 : rom_data = 10'b1101101111;
            10'd184 : rom_data = 10'b1101101111;
            10'd185 : rom_data = 10'b1100101111;
            10'd186 : rom_data = 10'b0100101101;
            10'd187 : rom_data = 10'b0100101101;
            10'd188 : rom_data = 10'b0100100001;
            10'd189 : rom_data = 10'b0000100000;
            10'd190 : rom_data = 10'b0000000000;
            10'd191 : rom_data = 10'b0000000000;
            10'd192 : rom_data = 10'b0000000000;
            10'd193 : rom_data = 10'b0000000000;
            10'd194 : rom_data = 10'b0000000000;
            10'd195 : rom_data = 10'b0000000000;
            10'd196 : rom_data = 10'b0000000000;
            10'd197 : rom_data = 10'b0000000000;
            10'd198 : rom_data = 10'b0000000000;
            10'd199 : rom_data = 10'b0000000000;
            10'd200 : rom_data = 10'b0000000000;
            10'd201 : rom_data = 10'b0000000000;
            10'd202 : rom_data = 10'b0000000000;
            10'd203 : rom_data = 10'b0000000000;
            10'd204 : rom_data = 10'b0000001000;
            10'd205 : rom_data = 10'b0000001100;
            10'd206 : rom_data = 10'b0100001101;
            10'd207 : rom_data = 10'b1110101101;
            10'd208 : rom_data = 10'b1111101101;
            10'd209 : rom_data = 10'b1111101101;
            10'd210 : rom_data = 10'b1111101111;
            10'd211 : rom_data = 10'b1111101111;
            10'd212 : rom_data = 10'b1110101111;
            10'd213 : rom_data = 10'b1110101111;
            10'd214 : rom_data = 10'b1110111101;
            10'd215 : rom_data = 10'b0100111101;
            10'd216 : rom_data = 10'b0100100001;
            10'd217 : rom_data = 10'b0000100001;
            10'd218 : rom_data = 10'b0000000000;
            10'd219 : rom_data = 10'b0000000000;
            10'd220 : rom_data = 10'b0000000000;
            10'd221 : rom_data = 10'b0000000000;
            10'd222 : rom_data = 10'b0000000000;
            10'd223 : rom_data = 10'b0000000000;
            10'd224 : rom_data = 10'b0000000000;
            10'd225 : rom_data = 10'b0000000000;
            10'd226 : rom_data = 10'b0000000000;
            10'd227 : rom_data = 10'b0000000000;
            10'd228 : rom_data = 10'b0000000000;
            10'd229 : rom_data = 10'b0000000000;
            10'd230 : rom_data = 10'b0000000000;
            10'd231 : rom_data = 10'b0000000000;
            10'd232 : rom_data = 10'b0010000000;
            10'd233 : rom_data = 10'b0010000000;
            10'd234 : rom_data = 10'b1110110001;
            10'd235 : rom_data = 10'b1111110101;
            10'd236 : rom_data = 10'b1111100001;
            10'd237 : rom_data = 10'b1111100001;
            10'd238 : rom_data = 10'b1111101011;
            10'd239 : rom_data = 10'b1110101111;
            10'd240 : rom_data = 10'b1110101111;
            10'd241 : rom_data = 10'b1110111111;
            10'd242 : rom_data = 10'b1110111101;
            10'd243 : rom_data = 10'b1110111101;
            10'd244 : rom_data = 10'b0110110001;
            10'd245 : rom_data = 10'b0100000001;
            10'd246 : rom_data = 10'b0000000000;
            10'd247 : rom_data = 10'b0000000000;
            10'd248 : rom_data = 10'b0000000000;
            10'd249 : rom_data = 10'b0000000000;
            10'd250 : rom_data = 10'b0000000000;
            10'd251 : rom_data = 10'b0000000000;
            10'd252 : rom_data = 10'b0000000000;
            10'd253 : rom_data = 10'b0000000000;
            10'd254 : rom_data = 10'b0000000000;
            10'd255 : rom_data = 10'b0000000000;
            10'd256 : rom_data = 10'b0000000000;
            10'd257 : rom_data = 10'b0000000000;
            10'd258 : rom_data = 10'b0000000000;
            10'd259 : rom_data = 10'b0010000000;
            10'd260 : rom_data = 10'b0010000000;
            10'd261 : rom_data = 10'b1110010001;
            10'd262 : rom_data = 10'b1111110001;
            10'd263 : rom_data = 10'b1111110001;
            10'd264 : rom_data = 10'b1111110001;
            10'd265 : rom_data = 10'b1111100001;
            10'd266 : rom_data = 10'b1011100011;
            10'd267 : rom_data = 10'b1010101011;
            10'd268 : rom_data = 10'b1010001111;
            10'd269 : rom_data = 10'b1110011111;
            10'd270 : rom_data = 10'b1110011101;
            10'd271 : rom_data = 10'b1110011101;
            10'd272 : rom_data = 10'b0110010001;
            10'd273 : rom_data = 10'b0100000001;
            10'd274 : rom_data = 10'b0000000001;
            10'd275 : rom_data = 10'b0000000000;
            10'd276 : rom_data = 10'b0000000000;
            10'd277 : rom_data = 10'b0000000000;
            10'd278 : rom_data = 10'b0000000000;
            10'd279 : rom_data = 10'b0000000000;
            10'd280 : rom_data = 10'b0000000000;
            10'd281 : rom_data = 10'b0000000000;
            10'd282 : rom_data = 10'b0000000000;
            10'd283 : rom_data = 10'b0000000000;
            10'd284 : rom_data = 10'b0000000000;
            10'd285 : rom_data = 10'b0000000000;
            10'd286 : rom_data = 10'b0000000000;
            10'd287 : rom_data = 10'b0010000000;
            10'd288 : rom_data = 10'b1010000001;
            10'd289 : rom_data = 10'b1110110001;
            10'd290 : rom_data = 10'b1111110001;
            10'd291 : rom_data = 10'b1111110001;
            10'd292 : rom_data = 10'b1111110001;
            10'd293 : rom_data = 10'b0011100011;
            10'd294 : rom_data = 10'b0010101011;
            10'd295 : rom_data = 10'b0010001010;
            10'd296 : rom_data = 10'b1010001110;
            10'd297 : rom_data = 10'b1110011110;
            10'd298 : rom_data = 10'b1110011101;
            10'd299 : rom_data = 10'b1110010101;
            10'd300 : rom_data = 10'b0110010001;
            10'd301 : rom_data = 10'b0000000001;
            10'd302 : rom_data = 10'b0000000001;
            10'd303 : rom_data = 10'b0000000000;
            10'd304 : rom_data = 10'b0000000000;
            10'd305 : rom_data = 10'b0000000000;
            10'd306 : rom_data = 10'b0000000000;
            10'd307 : rom_data = 10'b0000000000;
            10'd308 : rom_data = 10'b0000000000;
            10'd309 : rom_data = 10'b0000000000;
            10'd310 : rom_data = 10'b0000000000;
            10'd311 : rom_data = 10'b0000000000;
            10'd312 : rom_data = 10'b0000000000;
            10'd313 : rom_data = 10'b0000000000;
            10'd314 : rom_data = 10'b0000000000;
            10'd315 : rom_data = 10'b0000000000;
            10'd316 : rom_data = 10'b1010010001;
            10'd317 : rom_data = 10'b1111110001;
            10'd318 : rom_data = 10'b1111110001;
            10'd319 : rom_data = 10'b1101110001;
            10'd320 : rom_data = 10'b0101101001;
            10'd321 : rom_data = 10'b0101101010;
            10'd322 : rom_data = 10'b0000101010;
            10'd323 : rom_data = 10'b0000001010;
            10'd324 : rom_data = 10'b1110011110;
            10'd325 : rom_data = 10'b1110011100;
            10'd326 : rom_data = 10'b1110011100;
            10'd327 : rom_data = 10'b1110010101;
            10'd328 : rom_data = 10'b0110000001;
            10'd329 : rom_data = 10'b0000000001;
            10'd330 : rom_data = 10'b0000000001;
            10'd331 : rom_data = 10'b0000000000;
            10'd332 : rom_data = 10'b0000000000;
            10'd333 : rom_data = 10'b0000000000;
            10'd334 : rom_data = 10'b0000000000;
            10'd335 : rom_data = 10'b0000000000;
            10'd336 : rom_data = 10'b0000000000;
            10'd337 : rom_data = 10'b0000000000;
            10'd338 : rom_data = 10'b0000000000;
            10'd339 : rom_data = 10'b0000000000;
            10'd340 : rom_data = 10'b0000000000;
            10'd341 : rom_data = 10'b0000000000;
            10'd342 : rom_data = 10'b0000000000;
            10'd343 : rom_data = 10'b0000000001;
            10'd344 : rom_data = 10'b1000010001;
            10'd345 : rom_data = 10'b1001110001;
            10'd346 : rom_data = 10'b1101110001;
            10'd347 : rom_data = 10'b0101111001;
            10'd348 : rom_data = 10'b0101101000;
            10'd349 : rom_data = 10'b0100101010;
            10'd350 : rom_data = 10'b0100101010;
            10'd351 : rom_data = 10'b1100101010;
            10'd352 : rom_data = 10'b1110011110;
            10'd353 : rom_data = 10'b1111011100;
            10'd354 : rom_data = 10'b1111011100;
            10'd355 : rom_data = 10'b1111010101;
            10'd356 : rom_data = 10'b0000000001;
            10'd357 : rom_data = 10'b0000000001;
            10'd358 : rom_data = 10'b0000000001;
            10'd359 : rom_data = 10'b0000000001;
            10'd360 : rom_data = 10'b0000000000;
            10'd361 : rom_data = 10'b0000000000;
            10'd362 : rom_data = 10'b0000000000;
            10'd363 : rom_data = 10'b0000000000;
            10'd364 : rom_data = 10'b0000000000;
            10'd365 : rom_data = 10'b0000000000;
            10'd366 : rom_data = 10'b0000000000;
            10'd367 : rom_data = 10'b0000000000;
            10'd368 : rom_data = 10'b0000000000;
            10'd369 : rom_data = 10'b0000000000;
            10'd370 : rom_data = 10'b0000000000;
            10'd371 : rom_data = 10'b0000010001;
            10'd372 : rom_data = 10'b1001110001;
            10'd373 : rom_data = 10'b1001110001;
            10'd374 : rom_data = 10'b1101111001;
            10'd375 : rom_data = 10'b0101111001;
            10'd376 : rom_data = 10'b0101101000;
            10'd377 : rom_data = 10'b0100101010;
            10'd378 : rom_data = 10'b1100101010;
            10'd379 : rom_data = 10'b1101111110;
            10'd380 : rom_data = 10'b1111111110;
            10'd381 : rom_data = 10'b1111011100;
            10'd382 : rom_data = 10'b1111011100;
            10'd383 : rom_data = 10'b1011010101;
            10'd384 : rom_data = 10'b0001000001;
            10'd385 : rom_data = 10'b0000000001;
            10'd386 : rom_data = 10'b0000000001;
            10'd387 : rom_data = 10'b0000000001;
            10'd388 : rom_data = 10'b0000000000;
            10'd389 : rom_data = 10'b0000000000;
            10'd390 : rom_data = 10'b0000000000;
            10'd391 : rom_data = 10'b0000000000;
            10'd392 : rom_data = 10'b0000000000;
            10'd393 : rom_data = 10'b0000000000;
            10'd394 : rom_data = 10'b0000000000;
            10'd395 : rom_data = 10'b0000000000;
            10'd396 : rom_data = 10'b0000000000;
            10'd397 : rom_data = 10'b0000000000;
            10'd398 : rom_data = 10'b0000000001;
            10'd399 : rom_data = 10'b0000010001;
            10'd400 : rom_data = 10'b1001010001;
            10'd401 : rom_data = 10'b1001110001;
            10'd402 : rom_data = 10'b1101111001;
            10'd403 : rom_data = 10'b1101111000;
            10'd404 : rom_data = 10'b1101111000;
            10'd405 : rom_data = 10'b1101111110;
            10'd406 : rom_data = 10'b1101111110;
            10'd407 : rom_data = 10'b1111111110;
            10'd408 : rom_data = 10'b1111111100;
            10'd409 : rom_data = 10'b1111111100;
            10'd410 : rom_data = 10'b1011011100;
            10'd411 : rom_data = 10'b0011011001;
            10'd412 : rom_data = 10'b0001000001;
            10'd413 : rom_data = 10'b0001000001;
            10'd414 : rom_data = 10'b0000000001;
            10'd415 : rom_data = 10'b0000000000;
            10'd416 : rom_data = 10'b0000000000;
            10'd417 : rom_data = 10'b0000000000;
            10'd418 : rom_data = 10'b0000000000;
            10'd419 : rom_data = 10'b0000000000;
            10'd420 : rom_data = 10'b0000000000;
            10'd421 : rom_data = 10'b0000000000;
            10'd422 : rom_data = 10'b0000000000;
            10'd423 : rom_data = 10'b0000000000;
            10'd424 : rom_data = 10'b0000000000;
            10'd425 : rom_data = 10'b0000000000;
            10'd426 : rom_data = 10'b0000000001;
            10'd427 : rom_data = 10'b0000010001;
            10'd428 : rom_data = 10'b1001010001;
            10'd429 : rom_data = 10'b1001010001;
            10'd430 : rom_data = 10'b1001110100;
            10'd431 : rom_data = 10'b1101111100;
            10'd432 : rom_data = 10'b1101111110;
            10'd433 : rom_data = 10'b1101111110;
            10'd434 : rom_data = 10'b1101111110;
            10'd435 : rom_data = 10'b1111111110;
            10'd436 : rom_data = 10'b1111111100;
            10'd437 : rom_data = 10'b1111111100;
            10'd438 : rom_data = 10'b1011111100;
            10'd439 : rom_data = 10'b0001011001;
            10'd440 : rom_data = 10'b0001000001;
            10'd441 : rom_data = 10'b0001000001;
            10'd442 : rom_data = 10'b0000000001;
            10'd443 : rom_data = 10'b0000000000;
            10'd444 : rom_data = 10'b0000000000;
            10'd445 : rom_data = 10'b0000000000;
            10'd446 : rom_data = 10'b0000000000;
            10'd447 : rom_data = 10'b0000000000;
            10'd448 : rom_data = 10'b0000000000;
            10'd449 : rom_data = 10'b0000000000;
            10'd450 : rom_data = 10'b0000000000;
            10'd451 : rom_data = 10'b0000000000;
            10'd452 : rom_data = 10'b0000000000;
            10'd453 : rom_data = 10'b0000000000;
            10'd454 : rom_data = 10'b0000000001;
            10'd455 : rom_data = 10'b0000010001;
            10'd456 : rom_data = 10'b0001010101;
            10'd457 : rom_data = 10'b1001010101;
            10'd458 : rom_data = 10'b1101010100;
            10'd459 : rom_data = 10'b1101010100;
            10'd460 : rom_data = 10'b1101010110;
            10'd461 : rom_data = 10'b1101010110;
            10'd462 : rom_data = 10'b1111010110;
            10'd463 : rom_data = 10'b1111010110;
            10'd464 : rom_data = 10'b1111111100;
            10'd465 : rom_data = 10'b1111111100;
            10'd466 : rom_data = 10'b1011111101;
            10'd467 : rom_data = 10'b0001011001;
            10'd468 : rom_data = 10'b0001001001;
            10'd469 : rom_data = 10'b0001000001;
            10'd470 : rom_data = 10'b0000000001;
            10'd471 : rom_data = 10'b0000000000;
            10'd472 : rom_data = 10'b0000000000;
            10'd473 : rom_data = 10'b0000000000;
            10'd474 : rom_data = 10'b0000000000;
            10'd475 : rom_data = 10'b0000000000;
            10'd476 : rom_data = 10'b0000000000;
            10'd477 : rom_data = 10'b0000000000;
            10'd478 : rom_data = 10'b0000000000;
            10'd479 : rom_data = 10'b0000000000;
            10'd480 : rom_data = 10'b0000000000;
            10'd481 : rom_data = 10'b0000000001;
            10'd482 : rom_data = 10'b0000000001;
            10'd483 : rom_data = 10'b0000000101;
            10'd484 : rom_data = 10'b0001000101;
            10'd485 : rom_data = 10'b0001010101;
            10'd486 : rom_data = 10'b0101010100;
            10'd487 : rom_data = 10'b0101010100;
            10'd488 : rom_data = 10'b0101010110;
            10'd489 : rom_data = 10'b0101010110;
            10'd490 : rom_data = 10'b1111010110;
            10'd491 : rom_data = 10'b1111010110;
            10'd492 : rom_data = 10'b1111110100;
            10'd493 : rom_data = 10'b1111111101;
            10'd494 : rom_data = 10'b0001111101;
            10'd495 : rom_data = 10'b0001101101;
            10'd496 : rom_data = 10'b0001001001;
            10'd497 : rom_data = 10'b0001000001;
            10'd498 : rom_data = 10'b0000000000;
            10'd499 : rom_data = 10'b0000000000;
            10'd500 : rom_data = 10'b0000000000;
            10'd501 : rom_data = 10'b0000000000;
            10'd502 : rom_data = 10'b0000000000;
            10'd503 : rom_data = 10'b0000000000;
            10'd504 : rom_data = 10'b0000000000;
            10'd505 : rom_data = 10'b0000000000;
            10'd506 : rom_data = 10'b0000000000;
            10'd507 : rom_data = 10'b0000000000;
            10'd508 : rom_data = 10'b0000000000;
            10'd509 : rom_data = 10'b0000000001;
            10'd510 : rom_data = 10'b0000000101;
            10'd511 : rom_data = 10'b0000000101;
            10'd512 : rom_data = 10'b0001000101;
            10'd513 : rom_data = 10'b0101000101;
            10'd514 : rom_data = 10'b0101000100;
            10'd515 : rom_data = 10'b0101000110;
            10'd516 : rom_data = 10'b0101000110;
            10'd517 : rom_data = 10'b0111010110;
            10'd518 : rom_data = 10'b1111010110;
            10'd519 : rom_data = 10'b1111010110;
            10'd520 : rom_data = 10'b1111110101;
            10'd521 : rom_data = 10'b1111111101;
            10'd522 : rom_data = 10'b0001101101;
            10'd523 : rom_data = 10'b0001101101;
            10'd524 : rom_data = 10'b0001001101;
            10'd525 : rom_data = 10'b0000000001;
            10'd526 : rom_data = 10'b0000000000;
            10'd527 : rom_data = 10'b0000000000;
            10'd528 : rom_data = 10'b0000000000;
            10'd529 : rom_data = 10'b0000000000;
            10'd530 : rom_data = 10'b0000000000;
            10'd531 : rom_data = 10'b0000000000;
            10'd532 : rom_data = 10'b0000000000;
            10'd533 : rom_data = 10'b0000000000;
            10'd534 : rom_data = 10'b0000000000;
            10'd535 : rom_data = 10'b0000000000;
            10'd536 : rom_data = 10'b0000000000;
            10'd537 : rom_data = 10'b0000000000;
            10'd538 : rom_data = 10'b0000000101;
            10'd539 : rom_data = 10'b0000000101;
            10'd540 : rom_data = 10'b0101000101;
            10'd541 : rom_data = 10'b0101000101;
            10'd542 : rom_data = 10'b0101000101;
            10'd543 : rom_data = 10'b0101000110;
            10'd544 : rom_data = 10'b0101000110;
            10'd545 : rom_data = 10'b0011000110;
            10'd546 : rom_data = 10'b1011010110;
            10'd547 : rom_data = 10'b1111110101;
            10'd548 : rom_data = 10'b1111111101;
            10'd549 : rom_data = 10'b1101111101;
            10'd550 : rom_data = 10'b0001101101;
            10'd551 : rom_data = 10'b0001001101;
            10'd552 : rom_data = 10'b0001001101;
            10'd553 : rom_data = 10'b0000000100;
            10'd554 : rom_data = 10'b0000000000;
            10'd555 : rom_data = 10'b0000000000;
            10'd556 : rom_data = 10'b0000000000;
            10'd557 : rom_data = 10'b0000000000;
            10'd558 : rom_data = 10'b0000000000;
            10'd559 : rom_data = 10'b0000000000;
            10'd560 : rom_data = 10'b0000000000;
            10'd561 : rom_data = 10'b0000000000;
            10'd562 : rom_data = 10'b0000000000;
            10'd563 : rom_data = 10'b0000000000;
            10'd564 : rom_data = 10'b0000000000;
            10'd565 : rom_data = 10'b0000000000;
            10'd566 : rom_data = 10'b0000000101;
            10'd567 : rom_data = 10'b0000100101;
            10'd568 : rom_data = 10'b0100100101;
            10'd569 : rom_data = 10'b0101100101;
            10'd570 : rom_data = 10'b0101100101;
            10'd571 : rom_data = 10'b0101000111;
            10'd572 : rom_data = 10'b0111000111;
            10'd573 : rom_data = 10'b0011100111;
            10'd574 : rom_data = 10'b1111111111;
            10'd575 : rom_data = 10'b1111111101;
            10'd576 : rom_data = 10'b1111111101;
            10'd577 : rom_data = 10'b0101101101;
            10'd578 : rom_data = 10'b0001101101;
            10'd579 : rom_data = 10'b0000001101;
            10'd580 : rom_data = 10'b0000000100;
            10'd581 : rom_data = 10'b0000000000;
            10'd582 : rom_data = 10'b0000000000;
            10'd583 : rom_data = 10'b0000000000;
            10'd584 : rom_data = 10'b0000000000;
            10'd585 : rom_data = 10'b0000000000;
            10'd586 : rom_data = 10'b0000000000;
            10'd587 : rom_data = 10'b0000000000;
            10'd588 : rom_data = 10'b0000000000;
            10'd589 : rom_data = 10'b0000000000;
            10'd590 : rom_data = 10'b0000000000;
            10'd591 : rom_data = 10'b0000000000;
            10'd592 : rom_data = 10'b0000000000;
            10'd593 : rom_data = 10'b0000000000;
            10'd594 : rom_data = 10'b0000000001;
            10'd595 : rom_data = 10'b0000101101;
            10'd596 : rom_data = 10'b0100101101;
            10'd597 : rom_data = 10'b0100101101;
            10'd598 : rom_data = 10'b0101101111;
            10'd599 : rom_data = 10'b0101101111;
            10'd600 : rom_data = 10'b0111101111;
            10'd601 : rom_data = 10'b1111101111;
            10'd602 : rom_data = 10'b1111111111;
            10'd603 : rom_data = 10'b1111111101;
            10'd604 : rom_data = 10'b1101111101;
            10'd605 : rom_data = 10'b0101101101;
            10'd606 : rom_data = 10'b0000101101;
            10'd607 : rom_data = 10'b0000000100;
            10'd608 : rom_data = 10'b0000000000;
            10'd609 : rom_data = 10'b0000000000;
            10'd610 : rom_data = 10'b0000000000;
            10'd611 : rom_data = 10'b0000000000;
            10'd612 : rom_data = 10'b0000000000;
            10'd613 : rom_data = 10'b0000000000;
            10'd614 : rom_data = 10'b0000000000;
            10'd615 : rom_data = 10'b0000000000;
            10'd616 : rom_data = 10'b0000000000;
            10'd617 : rom_data = 10'b0000000000;
            10'd618 : rom_data = 10'b0000000000;
            10'd619 : rom_data = 10'b0000000000;
            10'd620 : rom_data = 10'b0000000000;
            10'd621 : rom_data = 10'b0000000000;
            10'd622 : rom_data = 10'b0000000000;
            10'd623 : rom_data = 10'b0000001001;
            10'd624 : rom_data = 10'b0100101101;
            10'd625 : rom_data = 10'b0100101101;
            10'd626 : rom_data = 10'b0100101111;
            10'd627 : rom_data = 10'b0110101111;
            10'd628 : rom_data = 10'b0110101111;
            10'd629 : rom_data = 10'b1110101011;
            10'd630 : rom_data = 10'b1110101011;
            10'd631 : rom_data = 10'b1110101001;
            10'd632 : rom_data = 10'b0100101001;
            10'd633 : rom_data = 10'b0100101001;
            10'd634 : rom_data = 10'b0000000000;
            10'd635 : rom_data = 10'b0000000000;
            10'd636 : rom_data = 10'b0000000000;
            10'd637 : rom_data = 10'b0000000000;
            10'd638 : rom_data = 10'b0000000000;
            10'd639 : rom_data = 10'b0000000000;
            10'd640 : rom_data = 10'b0000000000;
            10'd641 : rom_data = 10'b0000000000;
            10'd642 : rom_data = 10'b0000000000;
            10'd643 : rom_data = 10'b0000000000;
            10'd644 : rom_data = 10'b0000000000;
            10'd645 : rom_data = 10'b0000000000;
            10'd646 : rom_data = 10'b0000000000;
            10'd647 : rom_data = 10'b0000000000;
            10'd648 : rom_data = 10'b0000000000;
            10'd649 : rom_data = 10'b0000000000;
            10'd650 : rom_data = 10'b0000000000;
            10'd651 : rom_data = 10'b0000000000;
            10'd652 : rom_data = 10'b0000001000;
            10'd653 : rom_data = 10'b0100101001;
            10'd654 : rom_data = 10'b0100101001;
            10'd655 : rom_data = 10'b0110101001;
            10'd656 : rom_data = 10'b0110101001;
            10'd657 : rom_data = 10'b1110101001;
            10'd658 : rom_data = 10'b1110101001;
            10'd659 : rom_data = 10'b0100101001;
            10'd660 : rom_data = 10'b0100001000;
            10'd661 : rom_data = 10'b0000000000;
            10'd662 : rom_data = 10'b0000000000;
            10'd663 : rom_data = 10'b0000000000;
            10'd664 : rom_data = 10'b0000000000;
            10'd665 : rom_data = 10'b0000000000;
            10'd666 : rom_data = 10'b0000000000;
            10'd667 : rom_data = 10'b0000000000;
            10'd668 : rom_data = 10'b0000000000;
            10'd669 : rom_data = 10'b0000000000;
            10'd670 : rom_data = 10'b0000000000;
            10'd671 : rom_data = 10'b0000000000;
            10'd672 : rom_data = 10'b0000000000;
            10'd673 : rom_data = 10'b0000000000;
            10'd674 : rom_data = 10'b0000000000;
            10'd675 : rom_data = 10'b0000000000;
            10'd676 : rom_data = 10'b0000000000;
            10'd677 : rom_data = 10'b0000000000;
            10'd678 : rom_data = 10'b0000000000;
            10'd679 : rom_data = 10'b0000000000;
            10'd680 : rom_data = 10'b0000000000;
            10'd681 : rom_data = 10'b0000000000;
            10'd682 : rom_data = 10'b0000000000;
            10'd683 : rom_data = 10'b0110000000;
            10'd684 : rom_data = 10'b0110000000;
            10'd685 : rom_data = 10'b0110000000;
            10'd686 : rom_data = 10'b0100000000;
            10'd687 : rom_data = 10'b0000000000;
            10'd688 : rom_data = 10'b0000000000;
            10'd689 : rom_data = 10'b0000000000;
            10'd690 : rom_data = 10'b0000000000;
            10'd691 : rom_data = 10'b0000000000;
            10'd692 : rom_data = 10'b0000000000;
            10'd693 : rom_data = 10'b0000000000;
            10'd694 : rom_data = 10'b0000000000;
            10'd695 : rom_data = 10'b0000000000;
            10'd696 : rom_data = 10'b0000000000;
            10'd697 : rom_data = 10'b0000000000;
            10'd698 : rom_data = 10'b0000000000;
            10'd699 : rom_data = 10'b0000000000;
            10'd700 : rom_data = 10'b0000000000;
            10'd701 : rom_data = 10'b0000000000;
            10'd702 : rom_data = 10'b0000000000;
            10'd703 : rom_data = 10'b0000000000;
            10'd704 : rom_data = 10'b0000000000;
            10'd705 : rom_data = 10'b0000000000;
            10'd706 : rom_data = 10'b0000000000;
            10'd707 : rom_data = 10'b0000000000;
            10'd708 : rom_data = 10'b0000000000;
            10'd709 : rom_data = 10'b0000000000;
            10'd710 : rom_data = 10'b0000000000;
            10'd711 : rom_data = 10'b0000000000;
            10'd712 : rom_data = 10'b0000000000;
            10'd713 : rom_data = 10'b0000000000;
            10'd714 : rom_data = 10'b0000000000;
            10'd715 : rom_data = 10'b0000000000;
            10'd716 : rom_data = 10'b0000000000;
            10'd717 : rom_data = 10'b0000000000;
            10'd718 : rom_data = 10'b0000000000;
            10'd719 : rom_data = 10'b0000000000;
            10'd720 : rom_data = 10'b0000000000;
            10'd721 : rom_data = 10'b0000000000;
            10'd722 : rom_data = 10'b0000000000;
            10'd723 : rom_data = 10'b0000000000;
            10'd724 : rom_data = 10'b0000000000;
            10'd725 : rom_data = 10'b0000000000;
            10'd726 : rom_data = 10'b0000000000;
            10'd727 : rom_data = 10'b0000000000;
            10'd728 : rom_data = 10'b0000000000;
            10'd729 : rom_data = 10'b0000000000;
            10'd730 : rom_data = 10'b0000000000;
            10'd731 : rom_data = 10'b0000000000;
            10'd732 : rom_data = 10'b0000000000;
            10'd733 : rom_data = 10'b0000000000;
            10'd734 : rom_data = 10'b0000000000;
            10'd735 : rom_data = 10'b0000000000;
            10'd736 : rom_data = 10'b0000000000;
            10'd737 : rom_data = 10'b0000000000;
            10'd738 : rom_data = 10'b0000000000;
            10'd739 : rom_data = 10'b0000000000;
            10'd740 : rom_data = 10'b0000000000;
            10'd741 : rom_data = 10'b0000000000;
            10'd742 : rom_data = 10'b0000000000;
            10'd743 : rom_data = 10'b0000000000;
            10'd744 : rom_data = 10'b0000000000;
            10'd745 : rom_data = 10'b0000000000;
            10'd746 : rom_data = 10'b0000000000;
            10'd747 : rom_data = 10'b0000000000;
            10'd748 : rom_data = 10'b0000000000;
            10'd749 : rom_data = 10'b0000000000;
            10'd750 : rom_data = 10'b0000000000;
            10'd751 : rom_data = 10'b0000000000;
            10'd752 : rom_data = 10'b0000000000;
            10'd753 : rom_data = 10'b0000000000;
            10'd754 : rom_data = 10'b0000000000;
            10'd755 : rom_data = 10'b0000000000;
            10'd756 : rom_data = 10'b0000000000;
            10'd757 : rom_data = 10'b0000000000;
            10'd758 : rom_data = 10'b0000000000;
            10'd759 : rom_data = 10'b0000000000;
            10'd760 : rom_data = 10'b0000000000;
            10'd761 : rom_data = 10'b0000000000;
            10'd762 : rom_data = 10'b0000000000;
            10'd763 : rom_data = 10'b0000000000;
            10'd764 : rom_data = 10'b0000000000;
            10'd765 : rom_data = 10'b0000000000;
            10'd766 : rom_data = 10'b0000000000;
            10'd767 : rom_data = 10'b0000000000;
            10'd768 : rom_data = 10'b0000000000;
            10'd769 : rom_data = 10'b0000000000;
            10'd770 : rom_data = 10'b0000000000;
            10'd771 : rom_data = 10'b0000000000;
            10'd772 : rom_data = 10'b0000000000;
            10'd773 : rom_data = 10'b0000000000;
            10'd774 : rom_data = 10'b0000000000;
            10'd775 : rom_data = 10'b0000000000;
            10'd776 : rom_data = 10'b0000000000;
            10'd777 : rom_data = 10'b0000000000;
            10'd778 : rom_data = 10'b0000000000;
            10'd779 : rom_data = 10'b0000000000;
            10'd780 : rom_data = 10'b0000000000;
            10'd781 : rom_data = 10'b0000000000;
            10'd782 : rom_data = 10'b0000000000;
            10'd783 : rom_data = 10'b0000000000;
            default:  rom_data = 10'b0000000000;
        endcase
        end
    endfunction

    // Lógica de Visão Periférica (Borrar o molde para aceitar erros de alinhamento)
    always @(*) begin
        // Lê o centro
        rom_data = get_rom_data(ram_addr);
        
        // Lê a esquerda (cuidado com o zero)
        if (ram_addr > 0) 
            rom_data_left = get_rom_data(ram_addr - 10'd1);
        else 
            rom_data_left = 10'b0;
        
        // Lê a direita (cuidado com o 783)
        if (ram_addr < 783) 
            rom_data_right = get_rom_data(ram_addr + 10'd1);
        else 
            rom_data_right = 10'b0;
    end

    integer i;

    always @(posedge clk) begin
        if (!rst_n) begin
            state <= IDLE; ram_addr <= 0; prediction <= 0; done <= 0;
            total_ink <= 0;
            for (i=0; i<10; i=i+1) score[i] <= 0;
        end else begin
            case (state)
                IDLE: begin
                    done <= 0; ram_addr <= 0;
                    if (start) begin 
                        for (i=0; i<10; i=i+1) score[i] <= 0;
                        total_ink <= 0;
                        state <= WAIT_RAM;
                    end
                end

                WAIT_RAM: state <= CALC; 

                CALC: begin
                    // Se você desenhou TINTA (1)
                    if (ram_data == 1) begin
                        total_ink <= total_ink + 1;

                        for (i=0; i<10; i=i+1) begin
                            // TOLERÂNCIA ESPACIAL (O Segredo do Sucesso):
                            // Se o molde tiver tinta aqui, OU na esquerda, OU na direita, conta ponto.
                            // Isso faz o traço do "1" ficar mais grosso na memória da IA.
                            
                            if (rom_data[i] || rom_data_left[i] || rom_data_right[i]) begin
                                score[i] <= score[i] + 10; // ACERTOU!
                            end else begin
                                score[i] <= score[i] - 20; // ERROU! (Punição mais forte)
                            end
                        end
                    end 
                    // Se ram_data == 0, ignoramos.

                    if (ram_addr == 783) state <= RESULT;
                    else begin 
                        ram_addr <= ram_addr + 1;
                        state <= WAIT_RAM;
                    end
                end

                RESULT: begin
                    // Filtro de Ruído
                    if (total_ink < 5 || total_ink > 700) begin
                        prediction <= 15;
                    end else begin
                        prediction <= 0; 
                        if (score[1] >= score[0] && score[1] >= score[2] && score[1] >= score[3] && score[1] >= score[4] && score[1] >= score[5] && score[1] >= score[6] && score[1] >= score[7] && score[1] >= score[8] && score[1] >= score[9]) prediction <= 1;
                        else if (score[2] >= score[0] && score[2] >= score[3] && score[2] >= score[4] && score[2] >= score[5] && score[2] >= score[6] && score[2] >= score[7] && score[2] >= score[8] && score[2] >= score[9]) prediction <= 2;
                        else if (score[3] >= score[0] && score[3] >= score[4] && score[3] >= score[5] && score[3] >= score[6] && score[3] >= score[7] && score[3] >= score[8] && score[3] >= score[9]) prediction <= 3;
                        else if (score[4] >= score[0] && score[4] >= score[5] && score[4] >= score[6] && score[4] >= score[7] && score[4] >= score[8] && score[4] >= score[9]) prediction <= 4;
                        else if (score[5] >= score[0] && score[5] >= score[6] && score[5] >= score[7] && score[5] >= score[8] && score[5] >= score[9]) prediction <= 5;
                        else if (score[6] >= score[0] && score[6] >= score[7] && score[6] >= score[8] && score[6] >= score[9]) prediction <= 6;
                        else if (score[7] >= score[0] && score[7] >= score[8] && score[7] >= score[9]) prediction <= 7;
                        else if (score[8] >= score[0] && score[8] >= score[9]) prediction <= 8;
                        else if (score[9] >= score[0]) prediction <= 9;
                        else prediction <= 0;
                    end
                    
                    done <= 1; state <= IDLE;
                end
            endcase
        end
    end
endmodule